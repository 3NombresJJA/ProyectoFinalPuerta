library verilog;
use verilog.vl_types.all;
entity ProyectoFinal_vlg_vec_tst is
end ProyectoFinal_vlg_vec_tst;
