library verilog;
use verilog.vl_types.all;
entity ProyectoFinal_vlg_check_tst is
    port(
        Close           : in     vl_logic;
        Cont0           : in     vl_logic;
        Cont1           : in     vl_logic;
        Cont2           : in     vl_logic;
        Cont3           : in     vl_logic;
        \Open\          : in     vl_logic;
        Q0              : in     vl_logic;
        Q1              : in     vl_logic;
        Temp            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ProyectoFinal_vlg_check_tst;
